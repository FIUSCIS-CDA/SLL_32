//////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: MUX32_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbench();
`include "../Test/Test.v"

///////////////////////////////////////////////////////////////////////////////////
// Inputs: A (32 bits)
//         H (5 bits)
reg[31:0] A; 
reg[4:0] H;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Output: Y (32-bit)
wire[31:0] Y;
///////////////////////////////////////////////////////////////////////////////////

SLL_32 mySLL(.A(A),.H(H),.Y(Y));

initial begin

//////////////////////////////////////////////////////////////////////////////
// Initialize A
A = 47;
//////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////
//  Testing: All 5-bit S values 0 to 31
for (H=5'b00000; H <= 5'b11111; H = H + 5'b00001) begin
   $display("Testing: H=%b", H);
   #10;
   verifyEqual32(Y, A*(2**H));
   // You need this because the counter will reset to 0 otherwise
   if (H == 5'b11111) begin
    $display("All tests passed.");
    $stop;
   end
end
////////////////////////////////////////////////////////////////////////////////////////
  
end

endmodule